//created by zhouhang 20170216
//wave review 

module Wave_Review(
	clk_i,
	rst_n_i,
	
	rise_valid_i,
	fall_valid_i,
	gap_point_i,
	
	ask_o
);


endmodule
